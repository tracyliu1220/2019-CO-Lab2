module B_Control(
    zero_i,
    result_i,
    BranchType,
    control_o
);

//I/O ports
input         zero_i;
input  [31:0] result_i;
input         BranchType;
output        control_o;  

//Internal Signals

//Main function

endmodule